
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity cordic is
    Port (
        clk: in std_logic;
        rst: in std_logic
    );

end cordic;

architecture Behavioral of cordic is
begin
    
    process(clk)
    begin

    end process;
    
    
end Behavioral;
